Vim�UnDo� ���	t���4@�IϹ�J$`{�iK���J�G   	                 
       
   
   
    ^֚w    _�                             ����                                                                                                                                                                                                                                                                                                                                                             ^֙�     �                   5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             ^֙�     �                  module counter_165�_�                       "    ����                                                                                                                                                                                                                                                                                                                                                             ^֙�     �                  #module counter_16(clk, counter_out)5�_�                       #    ����                                                                                                                                                                                                                                                                                                                                                             ^֙�     �                  #module counter_16(clk, counter_out)5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             ^֙�     �                 output reg counter_out5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             ^֚@     �                 output reg counter_out[15:0]5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             ^֚A     �                 output reg counter_out[15:0]5�_�      	                     ����                                                                                                                                                                                                                                                                                                                                                             ^֚q     �                 always @5�_�      
           	          ����                                                                                                                                                                                                                                                                                                                                                             ^֚u     �                 always @(posedge clk)5�_�   	               
          ����                                                                                                                                                                                                                                                                                                                                                             ^֚v    �                 always @(posedge clk)5��